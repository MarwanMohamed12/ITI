module adder_4bit 
#(parameter n = 4)
(input clk,rst,
input [n-1:0]add1,
input [n-1:0]add2,
input carry_in,
output reg [n-1: 0] sum,
output reg carry_out
);
//-----------------------------







//write here combinational logic

//-----------------------------



always@(posedge clk)
begin
if(rst)begin

end

else
begin

end
end
endmodule
